.title KiCad schematic
.include "/media/fede/GIT/git/Simulacion-de-circuitos-electronicos/docs/KiCAD/library/LM741.MOD"
RL1 sal 0 10k
R3 Net-_R3-Pad1_ 0 3.9k
R2 sal Net-_R1-Pad1_ 100k
R1 Net-_R1-Pad1_ ent 4k
V3 ent 0 0 dc 0 ac 1 SIN(0 20m 1k)
V2 -Vcc 0 -15
V1 +Vcc 0 +15
XU1 Net-_R3-Pad1_ Net-_R1-Pad1_ +Vcc -Vcc sal LM741/NS
.ac dec 10 1 1MEG 
.end
